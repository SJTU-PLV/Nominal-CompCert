Require Import Coqlib Errors.
Require Import AST Linking Smallstep Invariant CallconvAlgebra.

Require Import Conventions Mach.
Require Import Locations.
Require Import LanguageInterface.

Require Import Integers.
Require Import Values Memory.

Require Import CallconvBig InjectFootprint Injp.
Require Import CAnew.
Require Import Asm Asmrel.
Require Import Asmgenproof0 Asmgenproof1.
Require Import Encrypt EncryptSpec Encryptproof.
Require Import Client Server.

Import GS.

(** 1st step : module linking *)
               
